`ifndef BP_ME_DEFINES_SVH
`define BP_ME_DEFINES_SVH

  `include "bsg_cache.vh"

  `include "bp_me_cce_defines.svh"
  `include "bp_me_cce_inst_defines.svh"
  `include "bp_me_cache_slice_defines.svh"

`endif

